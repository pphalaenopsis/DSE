LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY rangeComparator IS
PORT (
  NUM: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
  A: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
);
END rangeComparator;

ARCHITECTURE dataflow OF rangeComparator IS
BEGIN
  A(0) <= (NOT NUM(5) AND NOT NUM(4) AND NOT NUM(3)) OR 
        (NOT NUM(5) AND NOT NUM(4) AND NOT NUM(2) AND NOT NUM(1));
  A(1) <= (NOT NUM(5) AND NOT NUM(4) AND NUM(3) AND NUM(1)) OR
        (NOT NUM(5) AND NOT NUM(4) AND NUM(3) AND NUM(2)) OR
		  (NOT NUM(5) AND NUM(4) AND NOT NUM(3) AND NOT NUM(2));
		  
  A(2) <= (NOT NUM(5) AND NUM(4) AND NUM(3) AND NOT NUM(2)) OR
        (NOT NUM(5) AND NUM(4) AND NUM(2) AND NOT NUM(1)) OR
        (NOT NUM(5) AND NUM(4) AND NOT NUM(3) AND NUM(2));
  A(3) <= (NOT NUM(5) AND NUM(4) AND NUM(3) AND NUM(2) AND NUM(1)) OR
        (NUM(5) AND NOT NUM(4) AND NOT NUM(3));
  A(4) <= (NUM(5) AND NUM(4) AND NOT NUM(3) AND NOT NUM(2) AND NOT NUM(1)) OR
        (NUM(5) AND NOT NUM(4) AND NUM(3));
  A(5) <= (NUM(5) AND NUM(4) AND NOT NUM(3) AND NUM(2)) OR
        (NUM(5) AND NUM(4) AND NOT NUM(2) AND NUM(1)) OR
        (NUM(5) AND NUM(4) AND NUM(3)  AND NOT NUM(2));
  A(6) <= (NUM(5) AND NUM(4) AND NUM(3) AND NUM(2));

END dataflow;