LIBRARY ieee;
USE ieee.std_logic_1164.all;

-- "Empty" Entity
ENTITY Testbench_lab2_2 IS
END Testbench_lab2_2;

ARCHITECTURE Behavior OF Testbench_lab2_2 IS 

-- DUT
COMPONENT multi7seg
PORT (SW: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      HEX0,HEX1,HEX2,HEX3,HEX4: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END COMPONENT;

-- TESTBENCH SIGNALS
SIGNAL SEL_MUX: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL switches: STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL SEL_SHIFT: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL DISP0,DISP1,DISP2,DISP3,DISP4: STD_LOGIC_VECTOR(6 DOWNTO 0);

BEGIN 

PROCESS
BEGIN 
	SEL_MUX <= "00";
	SEL_SHIFT <= "000";
	WAIT FOR 20 ns;
	
	SEL_SHIFT <= "001";
	WAIT FOR 20 ns;
	
	SEL_SHIFT <= "010";
	WAIT FOR 20 ns;
	
	SEL_SHIFT <= "011";
	WAIT FOR 20 ns;
	
	SEL_SHIFT <= "100";
	WAIT;
END PROCESS;

switches <= SEL_SHIFT & SEL_MUX;

DECODER: multi7seg PORT MAP (switches,DISP0,DISP1,DISP2,DISP3,DISP4);

END Behavior;	