LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY BCD_converter is 
PORT ( SW: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
HEX0, HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END BCD_converter;

ARCHITECTURE Behavior OF BCD_converter IS


COMPONENT comparator IS
PORT(NUM: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
Z: OUT STD_LOGIC);
END COMPONENT;

COMPONENT circuit_A IS
PORT (DIGITS: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
A0,A1,A2: OUT STD_LOGIC);
END COMPONENT;

COMPONENT circuit_B IS
PORT (Z: IN STD_LOGIC;
DISPLAY: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END COMPONENT;

COMPONENT segment7 IS
PORT (M: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
DISPLAY: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END COMPONENT; 

COMPONENT mux IS
PORT (V,A : IN STD_LOGIC;
sel: IN STD_LOGIC;
M: OUT STD_LOGIC);
END COMPONENT; 

SIGNAL z: std_logic;
SIGNAL a0,a1,a2: std_logic;
SIGNAL m0,m1,m2,m3: std_logic;
SIGNAL digit: std_logic_vector(3 downto 0);

BEGIN 
COMP: comparator PORT MAP(SW(3 DOWNTO 0),z);
DISP1: circuit_B PORT MAP(z,HEX1(6 DOWNTO 0));
CIRA: circuit_A PORT MAP(SW(2 DOWNTO 0),a0,a1,a2);
MUX0: mux PORT MAP(SW(0),a0,z,m0);
MUX1: mux PORT MAP(SW(1),a1,z,m1);
MUX2: mux PORT MAP(SW(2),a2,z,m2);
MUX3: mux PORT MAP(SW(3),'0',z,m3);

digit <= m3 & m2 & m1 & m0;

DISP0: segment7 PORT MAP(digit,HEX0(6 DOWNTO 0));

END Behavior;